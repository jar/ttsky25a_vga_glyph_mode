VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO white_rabbit_small
  CLASS BLOCK ;
  FOREIGN white_rabbit_small ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.800 BY 14.280 ;
  OBS
      LAYER met1 ;
        RECT 0.000 14.000 3.640 14.280 ;
      LAYER met1 ;
        RECT 3.640 14.000 4.200 14.280 ;
      LAYER met1 ;
        RECT 0.000 13.720 3.360 14.000 ;
      LAYER met1 ;
        RECT 3.360 13.720 4.200 14.000 ;
      LAYER met1 ;
        RECT 0.000 13.160 3.080 13.720 ;
      LAYER met1 ;
        RECT 3.080 13.160 4.200 13.720 ;
      LAYER met1 ;
        RECT 4.200 13.440 9.800 14.280 ;
        RECT 4.200 13.160 5.880 13.440 ;
      LAYER met1 ;
        RECT 5.880 13.160 6.440 13.440 ;
      LAYER met1 ;
        RECT 0.000 12.600 2.800 13.160 ;
      LAYER met1 ;
        RECT 2.800 12.600 3.920 13.160 ;
      LAYER met1 ;
        RECT 3.920 12.880 5.320 13.160 ;
      LAYER met1 ;
        RECT 5.320 12.880 6.440 13.160 ;
      LAYER met1 ;
        RECT 6.440 12.880 9.800 13.440 ;
        RECT 3.920 12.600 4.760 12.880 ;
      LAYER met1 ;
        RECT 4.760 12.600 6.160 12.880 ;
      LAYER met1 ;
        RECT 6.160 12.600 9.800 12.880 ;
        RECT 0.000 11.200 2.520 12.600 ;
      LAYER met1 ;
        RECT 2.520 12.320 3.920 12.600 ;
      LAYER met1 ;
        RECT 3.920 12.320 4.480 12.600 ;
      LAYER met1 ;
        RECT 4.480 12.320 5.880 12.600 ;
        RECT 2.520 12.040 3.640 12.320 ;
      LAYER met1 ;
        RECT 3.640 12.040 4.200 12.320 ;
      LAYER met1 ;
        RECT 4.200 12.040 5.880 12.320 ;
      LAYER met1 ;
        RECT 5.880 12.040 9.800 12.600 ;
      LAYER met1 ;
        RECT 2.520 11.480 5.600 12.040 ;
      LAYER met1 ;
        RECT 5.600 11.480 9.800 12.040 ;
      LAYER met1 ;
        RECT 2.520 11.200 5.320 11.480 ;
      LAYER met1 ;
        RECT 5.320 11.200 9.800 11.480 ;
        RECT 0.000 10.920 2.240 11.200 ;
      LAYER met1 ;
        RECT 2.240 10.920 5.040 11.200 ;
      LAYER met1 ;
        RECT 5.040 10.920 9.800 11.200 ;
        RECT 0.000 10.640 1.400 10.920 ;
      LAYER met1 ;
        RECT 1.400 10.640 4.760 10.920 ;
      LAYER met1 ;
        RECT 4.760 10.640 9.800 10.920 ;
        RECT 0.000 10.360 1.120 10.640 ;
      LAYER met1 ;
        RECT 1.120 10.360 4.200 10.640 ;
      LAYER met1 ;
        RECT 0.000 10.080 0.840 10.360 ;
      LAYER met1 ;
        RECT 0.840 10.080 4.200 10.360 ;
      LAYER met1 ;
        RECT 0.000 9.800 0.560 10.080 ;
      LAYER met1 ;
        RECT 0.560 9.800 4.200 10.080 ;
      LAYER met1 ;
        RECT 0.000 9.520 0.280 9.800 ;
      LAYER met1 ;
        RECT 0.280 9.520 4.200 9.800 ;
        RECT 0.000 8.960 4.200 9.520 ;
      LAYER met1 ;
        RECT 0.000 8.400 0.280 8.960 ;
      LAYER met1 ;
        RECT 0.280 8.680 4.200 8.960 ;
      LAYER met1 ;
        RECT 4.200 8.680 9.800 10.640 ;
      LAYER met1 ;
        RECT 0.280 8.400 4.480 8.680 ;
      LAYER met1 ;
        RECT 4.480 8.400 9.800 8.680 ;
        RECT 0.000 8.120 0.560 8.400 ;
      LAYER met1 ;
        RECT 0.560 8.120 5.040 8.400 ;
      LAYER met1 ;
        RECT 5.040 8.120 9.800 8.400 ;
        RECT 0.000 6.440 1.400 8.120 ;
      LAYER met1 ;
        RECT 1.400 7.840 5.600 8.120 ;
      LAYER met1 ;
        RECT 5.600 7.840 9.800 8.120 ;
      LAYER met1 ;
        RECT 1.400 7.560 6.160 7.840 ;
      LAYER met1 ;
        RECT 6.160 7.560 9.800 7.840 ;
      LAYER met1 ;
        RECT 1.400 7.280 6.440 7.560 ;
      LAYER met1 ;
        RECT 6.440 7.280 9.800 7.560 ;
      LAYER met1 ;
        RECT 1.400 7.000 6.720 7.280 ;
      LAYER met1 ;
        RECT 6.720 7.000 9.800 7.280 ;
      LAYER met1 ;
        RECT 1.400 6.720 7.280 7.000 ;
      LAYER met1 ;
        RECT 7.280 6.720 9.800 7.000 ;
      LAYER met1 ;
        RECT 1.400 6.440 7.560 6.720 ;
      LAYER met1 ;
        RECT 7.560 6.440 9.800 6.720 ;
        RECT 0.000 5.040 1.120 6.440 ;
      LAYER met1 ;
        RECT 1.120 5.880 7.840 6.440 ;
      LAYER met1 ;
        RECT 7.840 5.880 9.800 6.440 ;
      LAYER met1 ;
        RECT 1.120 5.600 8.120 5.880 ;
      LAYER met1 ;
        RECT 8.120 5.600 9.800 5.880 ;
      LAYER met1 ;
        RECT 1.120 5.320 8.400 5.600 ;
      LAYER met1 ;
        RECT 8.400 5.320 9.800 5.600 ;
      LAYER met1 ;
        RECT 1.120 5.040 8.680 5.320 ;
      LAYER met1 ;
        RECT 0.000 4.200 1.400 5.040 ;
      LAYER met1 ;
        RECT 1.400 4.760 8.680 5.040 ;
      LAYER met1 ;
        RECT 8.680 4.760 9.800 5.320 ;
      LAYER met1 ;
        RECT 1.400 4.200 8.960 4.760 ;
      LAYER met1 ;
        RECT 0.000 3.920 1.680 4.200 ;
      LAYER met1 ;
        RECT 1.680 3.920 8.960 4.200 ;
      LAYER met1 ;
        RECT 8.960 3.920 9.800 4.760 ;
        RECT 0.000 1.120 1.960 3.920 ;
      LAYER met1 ;
        RECT 1.960 2.520 9.240 3.920 ;
      LAYER met1 ;
        RECT 9.240 2.520 9.800 3.920 ;
      LAYER met1 ;
        RECT 1.960 2.240 9.520 2.520 ;
      LAYER met1 ;
        RECT 9.520 2.240 9.800 2.520 ;
      LAYER met1 ;
        RECT 1.960 1.680 9.800 2.240 ;
        RECT 1.960 1.400 9.520 1.680 ;
      LAYER met1 ;
        RECT 9.520 1.400 9.800 1.680 ;
      LAYER met1 ;
        RECT 1.960 1.120 9.240 1.400 ;
      LAYER met1 ;
        RECT 0.000 0.560 1.400 1.120 ;
      LAYER met1 ;
        RECT 1.400 0.840 9.240 1.120 ;
      LAYER met1 ;
        RECT 9.240 0.840 9.800 1.400 ;
      LAYER met1 ;
        RECT 1.400 0.560 8.400 0.840 ;
      LAYER met1 ;
        RECT 8.400 0.560 9.800 0.840 ;
        RECT 0.000 0.280 1.120 0.560 ;
      LAYER met1 ;
        RECT 1.120 0.280 7.560 0.560 ;
      LAYER met1 ;
        RECT 7.560 0.280 9.800 0.560 ;
        RECT 0.000 0.000 1.400 0.280 ;
      LAYER met1 ;
        RECT 1.400 0.000 2.800 0.280 ;
      LAYER met1 ;
        RECT 2.800 0.000 3.080 0.280 ;
      LAYER met1 ;
        RECT 3.080 0.000 7.280 0.280 ;
      LAYER met1 ;
        RECT 7.280 0.000 9.800 0.280 ;
      LAYER met2 ;
        RECT 0.000 14.000 3.640 14.280 ;
      LAYER met2 ;
        RECT 3.640 14.000 4.200 14.280 ;
      LAYER met2 ;
        RECT 0.000 13.720 3.360 14.000 ;
      LAYER met2 ;
        RECT 3.360 13.720 4.200 14.000 ;
      LAYER met2 ;
        RECT 0.000 13.160 3.080 13.720 ;
      LAYER met2 ;
        RECT 3.080 13.160 4.200 13.720 ;
      LAYER met2 ;
        RECT 4.200 13.440 9.800 14.280 ;
        RECT 4.200 13.160 5.880 13.440 ;
      LAYER met2 ;
        RECT 5.880 13.160 6.440 13.440 ;
      LAYER met2 ;
        RECT 0.000 12.600 2.800 13.160 ;
      LAYER met2 ;
        RECT 2.800 12.600 3.920 13.160 ;
      LAYER met2 ;
        RECT 3.920 12.880 5.320 13.160 ;
      LAYER met2 ;
        RECT 5.320 12.880 6.440 13.160 ;
      LAYER met2 ;
        RECT 6.440 12.880 9.800 13.440 ;
        RECT 3.920 12.600 4.760 12.880 ;
      LAYER met2 ;
        RECT 4.760 12.600 6.160 12.880 ;
      LAYER met2 ;
        RECT 6.160 12.600 9.800 12.880 ;
        RECT 0.000 11.200 2.520 12.600 ;
      LAYER met2 ;
        RECT 2.520 12.320 3.920 12.600 ;
      LAYER met2 ;
        RECT 3.920 12.320 4.480 12.600 ;
      LAYER met2 ;
        RECT 4.480 12.320 5.880 12.600 ;
        RECT 2.520 12.040 3.640 12.320 ;
      LAYER met2 ;
        RECT 3.640 12.040 4.200 12.320 ;
      LAYER met2 ;
        RECT 4.200 12.040 5.880 12.320 ;
      LAYER met2 ;
        RECT 5.880 12.040 9.800 12.600 ;
      LAYER met2 ;
        RECT 2.520 11.480 5.600 12.040 ;
      LAYER met2 ;
        RECT 5.600 11.480 9.800 12.040 ;
      LAYER met2 ;
        RECT 2.520 11.200 5.320 11.480 ;
      LAYER met2 ;
        RECT 5.320 11.200 9.800 11.480 ;
        RECT 0.000 10.920 2.240 11.200 ;
      LAYER met2 ;
        RECT 2.240 10.920 5.040 11.200 ;
      LAYER met2 ;
        RECT 5.040 10.920 9.800 11.200 ;
        RECT 0.000 10.640 1.400 10.920 ;
      LAYER met2 ;
        RECT 1.400 10.640 4.760 10.920 ;
      LAYER met2 ;
        RECT 4.760 10.640 9.800 10.920 ;
        RECT 0.000 10.360 1.120 10.640 ;
      LAYER met2 ;
        RECT 1.120 10.360 4.200 10.640 ;
      LAYER met2 ;
        RECT 0.000 10.080 0.840 10.360 ;
      LAYER met2 ;
        RECT 0.840 10.080 4.200 10.360 ;
      LAYER met2 ;
        RECT 0.000 9.800 0.560 10.080 ;
      LAYER met2 ;
        RECT 0.560 9.800 4.200 10.080 ;
      LAYER met2 ;
        RECT 0.000 9.520 0.280 9.800 ;
      LAYER met2 ;
        RECT 0.280 9.520 4.200 9.800 ;
        RECT 0.000 8.960 4.200 9.520 ;
      LAYER met2 ;
        RECT 0.000 8.400 0.280 8.960 ;
      LAYER met2 ;
        RECT 0.280 8.680 4.200 8.960 ;
      LAYER met2 ;
        RECT 4.200 8.680 9.800 10.640 ;
      LAYER met2 ;
        RECT 0.280 8.400 4.480 8.680 ;
      LAYER met2 ;
        RECT 4.480 8.400 9.800 8.680 ;
        RECT 0.000 8.120 0.560 8.400 ;
      LAYER met2 ;
        RECT 0.560 8.120 5.040 8.400 ;
      LAYER met2 ;
        RECT 5.040 8.120 9.800 8.400 ;
        RECT 0.000 6.440 1.400 8.120 ;
      LAYER met2 ;
        RECT 1.400 7.840 5.600 8.120 ;
      LAYER met2 ;
        RECT 5.600 7.840 9.800 8.120 ;
      LAYER met2 ;
        RECT 1.400 7.560 6.160 7.840 ;
      LAYER met2 ;
        RECT 6.160 7.560 9.800 7.840 ;
      LAYER met2 ;
        RECT 1.400 7.280 6.440 7.560 ;
      LAYER met2 ;
        RECT 6.440 7.280 9.800 7.560 ;
      LAYER met2 ;
        RECT 1.400 7.000 6.720 7.280 ;
      LAYER met2 ;
        RECT 6.720 7.000 9.800 7.280 ;
      LAYER met2 ;
        RECT 1.400 6.720 7.280 7.000 ;
      LAYER met2 ;
        RECT 7.280 6.720 9.800 7.000 ;
      LAYER met2 ;
        RECT 1.400 6.440 7.560 6.720 ;
      LAYER met2 ;
        RECT 7.560 6.440 9.800 6.720 ;
        RECT 0.000 5.040 1.120 6.440 ;
      LAYER met2 ;
        RECT 1.120 5.880 7.840 6.440 ;
      LAYER met2 ;
        RECT 7.840 5.880 9.800 6.440 ;
      LAYER met2 ;
        RECT 1.120 5.600 8.120 5.880 ;
      LAYER met2 ;
        RECT 8.120 5.600 9.800 5.880 ;
      LAYER met2 ;
        RECT 1.120 5.320 8.400 5.600 ;
      LAYER met2 ;
        RECT 8.400 5.320 9.800 5.600 ;
      LAYER met2 ;
        RECT 1.120 5.040 8.680 5.320 ;
      LAYER met2 ;
        RECT 0.000 4.200 1.400 5.040 ;
      LAYER met2 ;
        RECT 1.400 4.760 8.680 5.040 ;
      LAYER met2 ;
        RECT 8.680 4.760 9.800 5.320 ;
      LAYER met2 ;
        RECT 1.400 4.200 8.960 4.760 ;
      LAYER met2 ;
        RECT 0.000 3.920 1.680 4.200 ;
      LAYER met2 ;
        RECT 1.680 3.920 8.960 4.200 ;
      LAYER met2 ;
        RECT 8.960 3.920 9.800 4.760 ;
        RECT 0.000 1.120 1.960 3.920 ;
      LAYER met2 ;
        RECT 1.960 2.520 9.240 3.920 ;
      LAYER met2 ;
        RECT 9.240 2.520 9.800 3.920 ;
      LAYER met2 ;
        RECT 1.960 2.240 9.520 2.520 ;
      LAYER met2 ;
        RECT 9.520 2.240 9.800 2.520 ;
      LAYER met2 ;
        RECT 1.960 1.680 9.800 2.240 ;
        RECT 1.960 1.400 9.520 1.680 ;
      LAYER met2 ;
        RECT 9.520 1.400 9.800 1.680 ;
      LAYER met2 ;
        RECT 1.960 1.120 9.240 1.400 ;
      LAYER met2 ;
        RECT 0.000 0.560 1.400 1.120 ;
      LAYER met2 ;
        RECT 1.400 0.840 9.240 1.120 ;
      LAYER met2 ;
        RECT 9.240 0.840 9.800 1.400 ;
      LAYER met2 ;
        RECT 1.400 0.560 8.400 0.840 ;
      LAYER met2 ;
        RECT 8.400 0.560 9.800 0.840 ;
        RECT 0.000 0.280 1.120 0.560 ;
      LAYER met2 ;
        RECT 1.120 0.280 7.560 0.560 ;
      LAYER met2 ;
        RECT 7.560 0.280 9.800 0.560 ;
        RECT 0.000 0.000 1.400 0.280 ;
      LAYER met2 ;
        RECT 1.400 0.000 2.800 0.280 ;
      LAYER met2 ;
        RECT 2.800 0.000 3.080 0.280 ;
      LAYER met2 ;
        RECT 3.080 0.000 7.280 0.280 ;
      LAYER met2 ;
        RECT 7.280 0.000 9.800 0.280 ;
      LAYER met3 ;
        RECT 0.000 0.000 9.800 14.280 ;
      LAYER met4 ;
        RECT 0.000 0.000 9.800 14.280 ;
      LAYER met5 ;
        RECT 0.000 0.000 9.800 14.280 ;
  END
END white_rabbit_small
END LIBRARY

