/*
 * Copyright (c) 2024 James Ross
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_vga_glyph_mode(
	input  wire [7:0] ui_in,    // Dedicated inputs
	output wire [7:0] uo_out,   // Dedicated outputs
	input  wire [7:0] uio_in,   // IOs: Input path
	output wire [7:0] uio_out,  // IOs: Output path
	output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
	input  wire       ena,      // always 1 when the design is powered, so you can ignore it
	input  wire       clk,      // clock
	input  wire       rst_n     // reset_n - low to reset
);

	// VGA signals
	wire hsync;
	wire vsync;
	wire [1:0] R;
	wire [1:0] G;
	wire [1:0] B;
	wire video_active;
	wire [9:0] pix_x;
	wire [9:0] pix_y;

	// TinyVGA PMOD
	assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

	// Unused outputs assigned to 0.
	assign uio_out = 0;
	assign uio_oe  = 0;

	wire [6:0] x_block = pix_x >> 3;
	wire [2:0] g_x = pix_x[2:0];
	wire [5:0] y_block = y_mem[pix_y >> 2];
	wire [3:0] g_y = pix_y - {y_block, 3'b000} - {1'b0, y_block, 2'b00};

	// Suppress unused signals warning
	wire _unused_ok = &{ena, ui_in, uio_in};

	reg [9:0] counter;

	hvsync_generator hvsync_gen(
		.clk(clk),
		.reset(~rst_n),
		.hsync(hsync),
		.vsync(vsync),
		.display_on(video_active),
		.hpos(pix_x),
		.vpos(pix_y)
	);
  
  wire [4:0] glyph_index = {x_block[2] ^ y_block[0]^counter[4], x_block[0] ^ y_block[1], x_block[1] ^ y_block[2], x_block[4] ^ y_block[3], x_block[3] ^ y_block[4]};
	  wire hl = g[glyph_index][g_y][g_x];
  wire [5:0] color = RGB[5];

	assign R = video_active ? {color[5] & hl, color[4] & hl} : 2'b00;
	assign G = video_active ? {color[3] & hl, color[2] & hl} : 2'b00;
	assign B = video_active ? {color[1] & hl, color[0] & hl} : 2'b00;
	
	always @(posedge vsync) begin
		if (~rst_n) begin
			counter <= 0;
		end else begin
			counter <= counter + 1;
		end
	end

  reg [5:0] RGB[0:7];
  initial begin
    RGB[0] = 6'b000000;
    RGB[1] = 6'b000100;
    RGB[2] = 6'b001000;
    RGB[3] = 6'b001100;
    RGB[4] = 6'b011100;
    RGB[5] = 6'b101101;
    RGB[6] = 6'b111110;
    RGB[7] = 6'b111111;
  end

	// glyphs
	reg [7:0] g[0:31][0:11];
	initial begin
    g[ 0][ 0] = 8'b00000000;
    g[ 0][ 1] = 8'b00011011;
    g[ 0][ 2] = 8'b00011011;
    g[ 0][ 3] = 8'b00011011;
    g[ 0][ 4] = 8'b00011011;
    g[ 0][ 5] = 8'b00110011;
    g[ 0][ 6] = 8'b00110011;
    g[ 0][ 7] = 8'b00110011;
    g[ 0][ 8] = 8'b01100001;
    g[ 0][ 9] = 8'b01100001;
    g[ 0][10] = 8'b01100001;
    g[ 0][11] = 8'b01100000;
    g[ 1][ 0] = 8'b00000000;
    g[ 1][ 1] = 8'b00000011;
    g[ 1][ 2] = 8'b00000011;
    g[ 1][ 3] = 8'b01111111;
    g[ 1][ 4] = 8'b01111111;
    g[ 1][ 5] = 8'b00000011;
    g[ 1][ 6] = 8'b00000011;
    g[ 1][ 7] = 8'b00000011;
    g[ 1][ 8] = 8'b00000011;
    g[ 1][ 9] = 8'b00000111;
    g[ 1][10] = 8'b01111110;
    g[ 1][11] = 8'b01111100;
    g[ 2][ 0] = 8'b00000000;
    g[ 2][ 1] = 8'b00001111;
    g[ 2][ 2] = 8'b00001111;
    g[ 2][ 3] = 8'b01000000;
    g[ 2][ 4] = 8'b01001111;
    g[ 2][ 5] = 8'b01001111;
    g[ 2][ 6] = 8'b01100000;
    g[ 2][ 7] = 8'b00100000;
    g[ 2][ 8] = 8'b00110000;
    g[ 2][ 9] = 8'b00111000;
    g[ 2][10] = 8'b00011111;
    g[ 2][11] = 8'b00001111;
    g[ 3][ 0] = 8'b00000000;
    g[ 3][ 1] = 8'b01100101;
    g[ 3][ 2] = 8'b01100101;
    g[ 3][ 3] = 8'b01101101;
    g[ 3][ 4] = 8'b01101011;
    g[ 3][ 5] = 8'b01101010;
    g[ 3][ 6] = 8'b01100000;
    g[ 3][ 7] = 8'b00110000;
    g[ 3][ 8] = 8'b00110000;
    g[ 3][ 9] = 8'b00110000;
    g[ 3][10] = 8'b00011000;
    g[ 3][11] = 8'b00011110;
    g[ 4][ 0] = 8'b00000000;
    g[ 4][ 1] = 8'b00001100;
    g[ 4][ 2] = 8'b00001100;
    g[ 4][ 3] = 8'b01111111;
    g[ 4][ 4] = 8'b01100011;
    g[ 4][ 5] = 8'b01100011;
    g[ 4][ 6] = 8'b01100000;
    g[ 4][ 7] = 8'b01100000;
    g[ 4][ 8] = 8'b01100000;
    g[ 4][ 9] = 8'b00110000;
    g[ 4][10] = 8'b00011000;
    g[ 4][11] = 8'b00001110;
    g[ 5][ 0] = 8'b00000000;
    g[ 5][ 1] = 8'b00011000;
    g[ 5][ 2] = 8'b00011000;
    g[ 5][ 3] = 8'b01111111;
    g[ 5][ 4] = 8'b01111111;
    g[ 5][ 5] = 8'b00011000;
    g[ 5][ 6] = 8'b00011000;
    g[ 5][ 7] = 8'b00011000;
    g[ 5][ 8] = 8'b00011100;
    g[ 5][ 9] = 8'b00001110;
    g[ 5][10] = 8'b00000011;
    g[ 5][11] = 8'b00000000;
    g[ 6][ 0] = 8'b00000000;
    g[ 6][ 1] = 8'b00000111;
    g[ 6][ 2] = 8'b00011100;
    g[ 6][ 3] = 8'b01110000;
    g[ 6][ 4] = 8'b00000000;
    g[ 6][ 5] = 8'b00000111;
    g[ 6][ 6] = 8'b00011100;
    g[ 6][ 7] = 8'b01110000;
    g[ 6][ 8] = 8'b00000000;
    g[ 6][ 9] = 8'b00000111;
    g[ 6][10] = 8'b00011100;
    g[ 6][11] = 8'b01110000;
    g[ 7][ 0] = 8'b00000000;
    g[ 7][ 1] = 8'b01111111;
    g[ 7][ 2] = 8'b00000110;
    g[ 7][ 3] = 8'b00000110;
    g[ 7][ 4] = 8'b01111111;
    g[ 7][ 5] = 8'b00000110;
    g[ 7][ 6] = 8'b00000110;
    g[ 7][ 7] = 8'b00000110;
    g[ 7][ 8] = 8'b00000110;
    g[ 7][ 9] = 8'b00001110;
    g[ 7][10] = 8'b01111100;
    g[ 7][11] = 8'b01111000;
    g[ 8][ 0] = 8'b00000000;
    g[ 8][ 1] = 8'b00000000;
    g[ 8][ 2] = 8'b00110110;
    g[ 8][ 3] = 8'b00110110;
    g[ 8][ 4] = 8'b01111111;
    g[ 8][ 5] = 8'b01111111;
    g[ 8][ 6] = 8'b00110110;
    g[ 8][ 7] = 8'b00110110;
    g[ 8][ 8] = 8'b00110000;
    g[ 8][ 9] = 8'b00110000;
    g[ 8][10] = 8'b00011000;
    g[ 8][11] = 8'b00001110;
    g[ 9][ 0] = 8'b00000000;
    g[ 9][ 1] = 8'b00000000;
    g[ 9][ 2] = 8'b01111111;
    g[ 9][ 3] = 8'b01100011;
    g[ 9][ 4] = 8'b01100011;
    g[ 9][ 5] = 8'b01100000;
    g[ 9][ 6] = 8'b01100000;
    g[ 9][ 7] = 8'b01100000;
    g[ 9][ 8] = 8'b01100000;
    g[ 9][ 9] = 8'b00110000;
    g[ 9][10] = 8'b00011000;
    g[ 9][11] = 8'b00001110;
    g[10][ 0] = 8'b00000000;
    g[10][ 1] = 8'b00110000;
    g[10][ 2] = 8'b00110000;
    g[10][ 3] = 8'b01111111;
    g[10][ 4] = 8'b01111111;
    g[10][ 5] = 8'b00110000;
    g[10][ 6] = 8'b00111000;
    g[10][ 7] = 8'b00111000;
    g[10][ 8] = 8'b00111100;
    g[10][ 9] = 8'b00110100;
    g[10][10] = 8'b00110110;
    g[10][11] = 8'b00110010;
    g[11][ 0] = 8'b00000000;
    g[11][ 1] = 8'b00000000;
    g[11][ 2] = 8'b01100011;
    g[11][ 3] = 8'b01100011;
    g[11][ 4] = 8'b01100011;
    g[11][ 5] = 8'b01100011;
    g[11][ 6] = 8'b01100011;
    g[11][ 7] = 8'b01100000;
    g[11][ 8] = 8'b01100000;
    g[11][ 9] = 8'b00110000;
    g[11][10] = 8'b00011000;
    g[11][11] = 8'b00001110;
    g[12][ 0] = 8'b00000000;
    g[12][ 1] = 8'b00001100;
    g[12][ 2] = 8'b01111111;
    g[12][ 3] = 8'b01111111;
    g[12][ 4] = 8'b00001100;
    g[12][ 5] = 8'b00001100;
    g[12][ 6] = 8'b00101101;
    g[12][ 7] = 8'b00101101;
    g[12][ 8] = 8'b00101101;
    g[12][ 9] = 8'b01101101;
    g[12][10] = 8'b01001101;
    g[12][11] = 8'b00011000;
    g[13][ 0] = 8'b00000000;
    g[13][ 1] = 8'b00000000;
    g[13][ 2] = 8'b01111110;
    g[13][ 3] = 8'b00111100;
    g[13][ 4] = 8'b01100000;
    g[13][ 5] = 8'b01100000;
    g[13][ 6] = 8'b01101100;
    g[13][ 7] = 8'b01101100;
    g[13][ 8] = 8'b00111100;
    g[13][ 9] = 8'b00011100;
    g[13][10] = 8'b00000110;
    g[13][11] = 8'b00000010;
    g[14][ 0] = 8'b00000000;
    g[14][ 1] = 8'b00000000;
    g[14][ 2] = 8'b00000110;
    g[14][ 3] = 8'b01111111;
    g[14][ 4] = 8'b01111111;
    g[14][ 5] = 8'b00001100;
    g[14][ 6] = 8'b00001100;
    g[14][ 7] = 8'b01111111;
    g[14][ 8] = 8'b01111111;
    g[14][ 9] = 8'b00011000;
    g[14][10] = 8'b00011000;
    g[14][11] = 8'b00011000;
    g[15][ 0] = 8'b00000000;
    g[15][ 1] = 8'b00000000;
    g[15][ 2] = 8'b00000000;
    g[15][ 3] = 8'b00001100;
    g[15][ 4] = 8'b00001100;
    g[15][ 5] = 8'b00001100;
    g[15][ 6] = 8'b00110110;
    g[15][ 7] = 8'b00110110;
    g[15][ 8] = 8'b01100110;
    g[15][ 9] = 8'b01110011;
    g[15][10] = 8'b01011011;
    g[15][11] = 8'b01001111;
    g[16][ 0] = 8'b00000000;
    g[16][ 1] = 8'b00000000;
    g[16][ 2] = 8'b01111110;
    g[16][ 3] = 8'b00000000;
    g[16][ 4] = 8'b00000000;
    g[16][ 5] = 8'b01111110;
    g[16][ 6] = 8'b00011000;
    g[16][ 7] = 8'b00011000;
    g[16][ 8] = 8'b00011000;
    g[16][ 9] = 8'b00011000;
    g[16][10] = 8'b00001100;
    g[16][11] = 8'b00000110;
    g[17][ 0] = 8'b00000000;
    g[17][ 1] = 8'b00001100;
    g[17][ 2] = 8'b00001100;
    g[17][ 3] = 8'b01111110;
    g[17][ 4] = 8'b01111110;
    g[17][ 5] = 8'b00011011;
    g[17][ 6] = 8'b00011001;
    g[17][ 7] = 8'b00011000;
    g[17][ 8] = 8'b00011000;
    g[17][ 9] = 8'b00011000;
    g[17][10] = 8'b00001100;
    g[17][11] = 8'b00000111;
    g[18][ 0] = 8'b00000000;
    g[18][ 1] = 8'b00000000;
    g[18][ 2] = 8'b00110000;
    g[18][ 3] = 8'b00110000;
    g[18][ 4] = 8'b00110010;
    g[18][ 5] = 8'b00110110;
    g[18][ 6] = 8'b00111100;
    g[18][ 7] = 8'b00111000;
    g[18][ 8] = 8'b01111000;
    g[18][ 9] = 8'b01011000;
    g[18][10] = 8'b00001100;
    g[18][11] = 8'b00000110;
    g[19][ 0] = 8'b00000000;
    g[19][ 1] = 8'b00000000;
    g[19][ 2] = 8'b00000110;
    g[19][ 3] = 8'b01111111;
    g[19][ 4] = 8'b01111111;
    g[19][ 5] = 8'b01100110;
    g[19][ 6] = 8'b01100110;
    g[19][ 7] = 8'b01100110;
    g[19][ 8] = 8'b01100110;
    g[19][ 9] = 8'b01100110;
    g[19][10] = 8'b01100010;
    g[19][11] = 8'b00111001;
    g[20][ 0] = 8'b00000000;
    g[20][ 1] = 8'b00000000;
    g[20][ 2] = 8'b01111110;
    g[20][ 3] = 8'b01111110;
    g[20][ 4] = 8'b00000000;
    g[20][ 5] = 8'b01111111;
    g[20][ 6] = 8'b01111111;
    g[20][ 7] = 8'b01100000;
    g[20][ 8] = 8'b01100000;
    g[20][ 9] = 8'b01110000;
    g[20][10] = 8'b00111000;
    g[20][11] = 8'b00011110;
    g[21][ 0] = 8'b00000000;
    g[21][ 1] = 8'b00000110;
    g[21][ 2] = 8'b00000110;
    g[21][ 3] = 8'b01111111;
    g[21][ 4] = 8'b01111111;
    g[21][ 5] = 8'b01100110;
    g[21][ 6] = 8'b01100110;
    g[21][ 7] = 8'b01100110;
    g[21][ 8] = 8'b00110110;
    g[21][ 9] = 8'b00000110;
    g[21][10] = 8'b01111110;
    g[21][11] = 8'b01111100;
    g[22][ 0] = 8'b00000000;
    g[22][ 1] = 8'b00001100;
    g[22][ 2] = 8'b01111111;
    g[22][ 3] = 8'b01111111;
    g[22][ 4] = 8'b01100000;
    g[22][ 5] = 8'b01100000;
    g[22][ 6] = 8'b01100000;
    g[22][ 7] = 8'b00110000;
    g[22][ 8] = 8'b00111100;
    g[22][ 9] = 8'b01101111;
    g[22][10] = 8'b01001100;
    g[22][11] = 8'b00001100;
    g[23][ 0] = 8'b00000000;
    g[23][ 1] = 8'b00000000;
    g[23][ 2] = 8'b00111110;
    g[23][ 3] = 8'b00111110;
    g[23][ 4] = 8'b00110000;
    g[23][ 5] = 8'b00110000;
    g[23][ 6] = 8'b00011000;
    g[23][ 7] = 8'b00011000;
    g[23][ 8] = 8'b00001100;
    g[23][ 9] = 8'b00011100;
    g[23][10] = 8'b00110110;
    g[23][11] = 8'b01100011;
    g[24][ 0] = 8'b00000000;
    g[24][ 1] = 8'b01111110;
    g[24][ 2] = 8'b01111110;
    g[24][ 3] = 8'b01100110;
    g[24][ 4] = 8'b01100011;
    g[24][ 5] = 8'b01100001;
    g[24][ 6] = 8'b01100100;
    g[24][ 7] = 8'b01111100;
    g[24][ 8] = 8'b00111000;
    g[24][ 9] = 8'b00011100;
    g[24][10] = 8'b00001110;
    g[24][11] = 8'b00000111;
    g[25][ 0] = 8'b00000000;
    g[25][ 1] = 8'b01111111;
    g[25][ 2] = 8'b01111111;
    g[25][ 3] = 8'b01100000;
    g[25][ 4] = 8'b01100000;
    g[25][ 5] = 8'b01100010;
    g[25][ 6] = 8'b01110110;
    g[25][ 7] = 8'b00111100;
    g[25][ 8] = 8'b00011000;
    g[25][ 9] = 8'b00111100;
    g[25][10] = 8'b01100110;
    g[25][11] = 8'b00000011;
    g[26][ 0] = 8'b00000000;
    g[26][ 1] = 8'b00111110;
    g[26][ 2] = 8'b01100011;
    g[26][ 3] = 8'b01100111;
    g[26][ 4] = 8'b01100111;
    g[26][ 5] = 8'b01101111;
    g[26][ 6] = 8'b01101011;
    g[26][ 7] = 8'b01111011;
    g[26][ 8] = 8'b01110011;
    g[26][ 9] = 8'b01110011;
    g[26][10] = 8'b01100011;
    g[26][11] = 8'b00111110;
    g[27][ 0] = 8'b00000000;
    g[27][ 1] = 8'b00001100;
    g[27][ 2] = 8'b00011100;
    g[27][ 3] = 8'b00011100;
    g[27][ 4] = 8'b00001100;
    g[27][ 5] = 8'b00001100;
    g[27][ 6] = 8'b00001100;
    g[27][ 7] = 8'b00001100;
    g[27][ 8] = 8'b00001100;
    g[27][ 9] = 8'b00001100;
    g[27][10] = 8'b00001100;
    g[27][11] = 8'b00001100;
    g[28][ 0] = 8'b00000000;
    g[28][ 1] = 8'b00111110;
    g[28][ 2] = 8'b01110001;
    g[28][ 3] = 8'b01100000;
    g[28][ 4] = 8'b01100000;
    g[28][ 5] = 8'b01100000;
    g[28][ 6] = 8'b00110000;
    g[28][ 7] = 8'b00011000;
    g[28][ 8] = 8'b00001100;
    g[28][ 9] = 8'b00000110;
    g[28][10] = 8'b00000011;
    g[28][11] = 8'b01111111;
    g[29][ 0] = 8'b00000000;
    g[29][ 1] = 8'b00111110;
    g[29][ 2] = 8'b01000011;
    g[29][ 3] = 8'b00000011;
    g[29][ 4] = 8'b00000011;
    g[29][ 5] = 8'b00000011;
    g[29][ 6] = 8'b00000110;
    g[29][ 7] = 8'b00011100;
    g[29][ 8] = 8'b00001100;
    g[29][ 9] = 8'b00000110;
    g[29][10] = 8'b00000011;
    g[29][11] = 8'b01111111;
    g[30][ 0] = 8'b00000000;
    g[30][ 1] = 8'b00000011;
    g[30][ 2] = 8'b00000111;
    g[30][ 3] = 8'b00001111;
    g[30][ 4] = 8'b00011011;
    g[30][ 5] = 8'b00110011;
    g[30][ 6] = 8'b01100011;
    g[30][ 7] = 8'b01100011;
    g[30][ 8] = 8'b01111111;
    g[30][ 9] = 8'b00000011;
    g[30][10] = 8'b00000011;
    g[30][11] = 8'b00000011;
    g[31][ 0] = 8'b00000000;
    g[31][ 1] = 8'b01111111;
    g[31][ 2] = 8'b00000011;
    g[31][ 3] = 8'b00000011;
    g[31][ 4] = 8'b00011111;
    g[31][ 5] = 8'b00111111;
    g[31][ 6] = 8'b01110000;
    g[31][ 7] = 8'b01100000;
    g[31][ 8] = 8'b01100000;
    g[31][ 9] = 8'b01100000;
    g[31][10] = 8'b01100001;
    g[31][11] = 8'b00111110;
	end

	// Division-by-3 lookup
	reg [5:0] y_mem[0:119];
	initial begin
		y_mem[0] = 6'd0;
		y_mem[1] = 6'd0;
		y_mem[2] = 6'd0;
		y_mem[3] = 6'd1;
		y_mem[4] = 6'd1;
		y_mem[5] = 6'd1;
		y_mem[6] = 6'd2;
		y_mem[7] = 6'd2;
		y_mem[8] = 6'd2;
		y_mem[9] = 6'd3;
		y_mem[10] = 6'd3;
		y_mem[11] = 6'd3;
		y_mem[12] = 6'd4;
		y_mem[13] = 6'd4;
		y_mem[14] = 6'd4;
		y_mem[15] = 6'd5;
		y_mem[16] = 6'd5;
		y_mem[17] = 6'd5;
		y_mem[18] = 6'd6;
		y_mem[19] = 6'd6;
		y_mem[20] = 6'd6;
		y_mem[21] = 6'd7;
		y_mem[22] = 6'd7;
		y_mem[23] = 6'd7;
		y_mem[24] = 6'd8;
		y_mem[25] = 6'd8;
		y_mem[26] = 6'd8;
		y_mem[27] = 6'd9;
		y_mem[28] = 6'd9;
		y_mem[29] = 6'd9;
		y_mem[30] = 6'd10;
		y_mem[31] = 6'd10;
		y_mem[32] = 6'd10;
		y_mem[33] = 6'd11;
		y_mem[34] = 6'd11;
		y_mem[35] = 6'd11;
		y_mem[36] = 6'd12;
		y_mem[37] = 6'd12;
		y_mem[38] = 6'd12;
		y_mem[39] = 6'd13;
		y_mem[40] = 6'd13;
		y_mem[41] = 6'd13;
		y_mem[42] = 6'd14;
		y_mem[43] = 6'd14;
		y_mem[44] = 6'd14;
		y_mem[45] = 6'd15;
		y_mem[46] = 6'd15;
		y_mem[47] = 6'd15;
		y_mem[48] = 6'd16;
		y_mem[49] = 6'd16;
		y_mem[50] = 6'd16;
		y_mem[51] = 6'd17;
		y_mem[52] = 6'd17;
		y_mem[53] = 6'd17;
		y_mem[54] = 6'd18;
		y_mem[55] = 6'd18;
		y_mem[56] = 6'd18;
		y_mem[57] = 6'd19;
		y_mem[58] = 6'd19;
		y_mem[59] = 6'd19;
		y_mem[60] = 6'd20;
		y_mem[61] = 6'd20;
		y_mem[62] = 6'd20;
		y_mem[63] = 6'd21;
		y_mem[64] = 6'd21;
		y_mem[65] = 6'd21;
		y_mem[66] = 6'd22;
		y_mem[67] = 6'd22;
		y_mem[68] = 6'd22;
		y_mem[69] = 6'd23;
		y_mem[70] = 6'd23;
		y_mem[71] = 6'd23;
		y_mem[72] = 6'd24;
		y_mem[73] = 6'd24;
		y_mem[74] = 6'd24;
		y_mem[75] = 6'd25;
		y_mem[76] = 6'd25;
		y_mem[77] = 6'd25;
		y_mem[78] = 6'd26;
		y_mem[79] = 6'd26;
		y_mem[80] = 6'd26;
		y_mem[81] = 6'd27;
		y_mem[82] = 6'd27;
		y_mem[83] = 6'd27;
		y_mem[84] = 6'd28;
		y_mem[85] = 6'd28;
		y_mem[86] = 6'd28;
		y_mem[87] = 6'd29;
		y_mem[88] = 6'd29;
		y_mem[89] = 6'd29;
		y_mem[90] = 6'd30;
		y_mem[91] = 6'd30;
		y_mem[92] = 6'd30;
		y_mem[93] = 6'd31;
		y_mem[94] = 6'd31;
		y_mem[95] = 6'd31;
		y_mem[96] = 6'd32;
		y_mem[97] = 6'd32;
		y_mem[98] = 6'd32;
		y_mem[99] = 6'd33;
		y_mem[100] = 6'd33;
		y_mem[101] = 6'd33;
		y_mem[102] = 6'd34;
		y_mem[103] = 6'd34;
		y_mem[104] = 6'd34;
		y_mem[105] = 6'd35;
		y_mem[106] = 6'd35;
		y_mem[107] = 6'd35;
		y_mem[108] = 6'd36;
		y_mem[109] = 6'd36;
		y_mem[110] = 6'd36;
		y_mem[111] = 6'd37;
		y_mem[112] = 6'd37;
		y_mem[113] = 6'd37;
		y_mem[114] = 6'd38;
		y_mem[115] = 6'd38;
		y_mem[116] = 6'd38;
		y_mem[117] = 6'd39;
		y_mem[118] = 6'd39;
		y_mem[119] = 6'd39;
	end

endmodule
