VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO white_rabbit
  CLASS BLOCK ;
  FOREIGN white_rabbit ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.760 BY 27.720 ;
  OBS
      LAYER met1 ;
        RECT 0.000 27.440 7.560 27.720 ;
      LAYER met1 ;
        RECT 7.560 27.440 8.120 27.720 ;
      LAYER met1 ;
        RECT 0.000 27.160 7.000 27.440 ;
      LAYER met1 ;
        RECT 7.000 27.160 8.120 27.440 ;
      LAYER met1 ;
        RECT 0.000 26.880 6.720 27.160 ;
      LAYER met1 ;
        RECT 6.720 26.880 8.120 27.160 ;
      LAYER met1 ;
        RECT 0.000 26.600 6.440 26.880 ;
      LAYER met1 ;
        RECT 6.440 26.600 8.120 26.880 ;
      LAYER met1 ;
        RECT 0.000 26.320 6.160 26.600 ;
      LAYER met1 ;
        RECT 6.160 26.320 8.120 26.600 ;
      LAYER met1 ;
        RECT 0.000 26.040 5.880 26.320 ;
      LAYER met1 ;
        RECT 5.880 26.040 8.120 26.320 ;
      LAYER met1 ;
        RECT 8.120 26.040 18.760 27.720 ;
        RECT 0.000 25.480 5.600 26.040 ;
      LAYER met1 ;
        RECT 5.600 25.480 8.120 26.040 ;
      LAYER met1 ;
        RECT 8.120 25.760 11.480 26.040 ;
      LAYER met1 ;
        RECT 11.480 25.760 12.040 26.040 ;
      LAYER met1 ;
        RECT 8.120 25.480 10.920 25.760 ;
      LAYER met1 ;
        RECT 10.920 25.480 12.040 25.760 ;
      LAYER met1 ;
        RECT 0.000 24.920 5.320 25.480 ;
      LAYER met1 ;
        RECT 5.320 24.920 7.840 25.480 ;
      LAYER met1 ;
        RECT 7.840 25.200 10.080 25.480 ;
      LAYER met1 ;
        RECT 10.080 25.200 12.040 25.480 ;
      LAYER met1 ;
        RECT 7.840 24.920 9.800 25.200 ;
      LAYER met1 ;
        RECT 9.800 24.920 12.040 25.200 ;
      LAYER met1 ;
        RECT 12.040 24.920 18.760 26.040 ;
        RECT 0.000 24.080 5.040 24.920 ;
      LAYER met1 ;
        RECT 5.040 24.640 7.840 24.920 ;
      LAYER met1 ;
        RECT 7.840 24.640 9.240 24.920 ;
      LAYER met1 ;
        RECT 9.240 24.640 11.760 24.920 ;
        RECT 5.040 24.080 7.560 24.640 ;
      LAYER met1 ;
        RECT 7.560 24.360 8.960 24.640 ;
      LAYER met1 ;
        RECT 8.960 24.360 11.760 24.640 ;
      LAYER met1 ;
        RECT 7.560 24.080 8.400 24.360 ;
      LAYER met1 ;
        RECT 8.400 24.080 11.760 24.360 ;
      LAYER met1 ;
        RECT 11.760 24.080 18.760 24.920 ;
        RECT 0.000 21.560 4.760 24.080 ;
      LAYER met1 ;
        RECT 4.760 23.800 7.560 24.080 ;
      LAYER met1 ;
        RECT 7.560 23.800 8.120 24.080 ;
      LAYER met1 ;
        RECT 8.120 23.800 11.480 24.080 ;
        RECT 4.760 23.240 7.280 23.800 ;
      LAYER met1 ;
        RECT 7.280 23.520 7.840 23.800 ;
      LAYER met1 ;
        RECT 7.840 23.520 11.480 23.800 ;
      LAYER met1 ;
        RECT 11.480 23.520 18.760 24.080 ;
        RECT 7.280 23.240 7.560 23.520 ;
      LAYER met1 ;
        RECT 7.560 23.240 11.200 23.520 ;
        RECT 4.760 22.960 11.200 23.240 ;
      LAYER met1 ;
        RECT 11.200 22.960 18.760 23.520 ;
      LAYER met1 ;
        RECT 4.760 22.680 10.920 22.960 ;
      LAYER met1 ;
        RECT 10.920 22.680 18.760 22.960 ;
      LAYER met1 ;
        RECT 4.760 22.120 10.640 22.680 ;
      LAYER met1 ;
        RECT 10.640 22.120 18.760 22.680 ;
      LAYER met1 ;
        RECT 4.760 21.840 10.360 22.120 ;
      LAYER met1 ;
        RECT 10.360 21.840 18.760 22.120 ;
      LAYER met1 ;
        RECT 4.760 21.560 10.080 21.840 ;
      LAYER met1 ;
        RECT 10.080 21.560 18.760 21.840 ;
        RECT 0.000 21.280 3.920 21.560 ;
      LAYER met1 ;
        RECT 3.920 21.280 9.800 21.560 ;
      LAYER met1 ;
        RECT 9.800 21.280 18.760 21.560 ;
        RECT 0.000 21.000 3.080 21.280 ;
      LAYER met1 ;
        RECT 3.080 21.000 9.520 21.280 ;
      LAYER met1 ;
        RECT 9.520 21.000 18.760 21.280 ;
        RECT 0.000 20.720 2.800 21.000 ;
      LAYER met1 ;
        RECT 2.800 20.720 8.960 21.000 ;
      LAYER met1 ;
        RECT 8.960 20.720 18.760 21.000 ;
        RECT 0.000 20.440 2.240 20.720 ;
      LAYER met1 ;
        RECT 2.240 20.440 8.680 20.720 ;
      LAYER met1 ;
        RECT 8.680 20.440 18.760 20.720 ;
        RECT 0.000 20.160 1.960 20.440 ;
      LAYER met1 ;
        RECT 1.960 20.160 8.120 20.440 ;
      LAYER met1 ;
        RECT 0.000 19.880 1.680 20.160 ;
      LAYER met1 ;
        RECT 1.680 19.880 8.120 20.160 ;
      LAYER met1 ;
        RECT 0.000 19.600 1.400 19.880 ;
      LAYER met1 ;
        RECT 1.400 19.600 8.120 19.880 ;
      LAYER met1 ;
        RECT 8.120 19.600 18.760 20.440 ;
        RECT 0.000 19.320 1.120 19.600 ;
      LAYER met1 ;
        RECT 1.120 19.320 8.400 19.600 ;
      LAYER met1 ;
        RECT 0.000 19.040 0.840 19.320 ;
      LAYER met1 ;
        RECT 0.840 19.040 8.400 19.320 ;
      LAYER met1 ;
        RECT 0.000 18.760 0.560 19.040 ;
      LAYER met1 ;
        RECT 0.560 18.760 8.400 19.040 ;
      LAYER met1 ;
        RECT 0.000 18.480 0.280 18.760 ;
      LAYER met1 ;
        RECT 0.280 18.480 8.400 18.760 ;
        RECT 0.000 17.360 8.400 18.480 ;
      LAYER met1 ;
        RECT 0.000 16.800 0.280 17.360 ;
      LAYER met1 ;
        RECT 0.280 16.800 8.400 17.360 ;
      LAYER met1 ;
        RECT 8.400 16.800 18.760 19.600 ;
        RECT 0.000 16.240 0.560 16.800 ;
      LAYER met1 ;
        RECT 0.560 16.520 8.680 16.800 ;
      LAYER met1 ;
        RECT 8.680 16.520 18.760 16.800 ;
      LAYER met1 ;
        RECT 0.560 16.240 9.240 16.520 ;
      LAYER met1 ;
        RECT 9.240 16.240 18.760 16.520 ;
        RECT 0.000 15.960 0.840 16.240 ;
      LAYER met1 ;
        RECT 0.840 15.960 9.800 16.240 ;
      LAYER met1 ;
        RECT 9.800 15.960 18.760 16.240 ;
        RECT 0.000 15.680 1.400 15.960 ;
      LAYER met1 ;
        RECT 1.400 15.680 10.360 15.960 ;
      LAYER met1 ;
        RECT 10.360 15.680 18.760 15.960 ;
        RECT 0.000 14.280 2.520 15.680 ;
      LAYER met1 ;
        RECT 2.520 15.400 10.920 15.680 ;
      LAYER met1 ;
        RECT 10.920 15.400 18.760 15.680 ;
      LAYER met1 ;
        RECT 2.520 15.120 11.200 15.400 ;
      LAYER met1 ;
        RECT 11.200 15.120 18.760 15.400 ;
      LAYER met1 ;
        RECT 2.520 14.840 11.760 15.120 ;
      LAYER met1 ;
        RECT 11.760 14.840 18.760 15.120 ;
      LAYER met1 ;
        RECT 2.520 14.560 12.040 14.840 ;
      LAYER met1 ;
        RECT 12.040 14.560 18.760 14.840 ;
      LAYER met1 ;
        RECT 2.520 14.280 12.600 14.560 ;
      LAYER met1 ;
        RECT 12.600 14.280 18.760 14.560 ;
        RECT 0.000 9.240 2.240 14.280 ;
      LAYER met1 ;
        RECT 2.240 14.000 12.880 14.280 ;
      LAYER met1 ;
        RECT 12.880 14.000 18.760 14.280 ;
      LAYER met1 ;
        RECT 2.240 13.720 13.160 14.000 ;
      LAYER met1 ;
        RECT 13.160 13.720 18.760 14.000 ;
      LAYER met1 ;
        RECT 2.240 13.440 13.440 13.720 ;
      LAYER met1 ;
        RECT 13.440 13.440 18.760 13.720 ;
      LAYER met1 ;
        RECT 2.240 13.160 13.720 13.440 ;
      LAYER met1 ;
        RECT 13.720 13.160 18.760 13.440 ;
      LAYER met1 ;
        RECT 2.240 12.880 14.000 13.160 ;
      LAYER met1 ;
        RECT 14.000 12.880 18.760 13.160 ;
      LAYER met1 ;
        RECT 2.240 12.600 14.280 12.880 ;
      LAYER met1 ;
        RECT 14.280 12.600 18.760 12.880 ;
      LAYER met1 ;
        RECT 2.240 12.320 14.560 12.600 ;
      LAYER met1 ;
        RECT 14.560 12.320 18.760 12.600 ;
      LAYER met1 ;
        RECT 2.240 12.040 14.840 12.320 ;
      LAYER met1 ;
        RECT 14.840 12.040 18.760 12.320 ;
      LAYER met1 ;
        RECT 2.240 11.760 15.120 12.040 ;
      LAYER met1 ;
        RECT 15.120 11.760 18.760 12.040 ;
      LAYER met1 ;
        RECT 2.240 11.480 15.400 11.760 ;
      LAYER met1 ;
        RECT 15.400 11.480 18.760 11.760 ;
      LAYER met1 ;
        RECT 2.240 11.200 15.680 11.480 ;
      LAYER met1 ;
        RECT 15.680 11.200 18.760 11.480 ;
      LAYER met1 ;
        RECT 2.240 10.640 15.960 11.200 ;
      LAYER met1 ;
        RECT 15.960 10.640 18.760 11.200 ;
      LAYER met1 ;
        RECT 2.240 10.360 16.240 10.640 ;
      LAYER met1 ;
        RECT 16.240 10.360 18.760 10.640 ;
      LAYER met1 ;
        RECT 2.240 9.800 16.520 10.360 ;
      LAYER met1 ;
        RECT 16.520 9.800 18.760 10.360 ;
      LAYER met1 ;
        RECT 2.240 9.240 16.800 9.800 ;
      LAYER met1 ;
        RECT 16.800 9.240 18.760 9.800 ;
        RECT 0.000 8.400 2.520 9.240 ;
      LAYER met1 ;
        RECT 2.520 8.680 17.080 9.240 ;
      LAYER met1 ;
        RECT 17.080 8.680 18.760 9.240 ;
      LAYER met1 ;
        RECT 2.520 8.400 17.360 8.680 ;
      LAYER met1 ;
        RECT 0.000 7.840 2.800 8.400 ;
      LAYER met1 ;
        RECT 2.800 8.120 17.360 8.400 ;
      LAYER met1 ;
        RECT 17.360 8.120 18.760 8.680 ;
      LAYER met1 ;
        RECT 2.800 7.840 17.640 8.120 ;
      LAYER met1 ;
        RECT 0.000 3.920 3.360 7.840 ;
      LAYER met1 ;
        RECT 3.360 7.000 17.640 7.840 ;
      LAYER met1 ;
        RECT 17.640 7.000 18.760 8.120 ;
      LAYER met1 ;
        RECT 3.360 4.200 17.920 7.000 ;
      LAYER met1 ;
        RECT 17.920 4.200 18.760 7.000 ;
      LAYER met1 ;
        RECT 3.360 3.920 18.480 4.200 ;
      LAYER met1 ;
        RECT 18.480 3.920 18.760 4.200 ;
        RECT 0.000 2.240 3.640 3.920 ;
      LAYER met1 ;
        RECT 3.640 3.080 18.760 3.920 ;
        RECT 3.640 2.800 18.480 3.080 ;
      LAYER met1 ;
        RECT 18.480 2.800 18.760 3.080 ;
      LAYER met1 ;
        RECT 3.640 2.240 17.920 2.800 ;
      LAYER met1 ;
        RECT 17.920 2.240 18.760 2.800 ;
        RECT 0.000 1.960 2.800 2.240 ;
      LAYER met1 ;
        RECT 2.800 1.960 17.640 2.240 ;
      LAYER met1 ;
        RECT 17.640 1.960 18.760 2.240 ;
        RECT 0.000 1.680 2.520 1.960 ;
      LAYER met1 ;
        RECT 2.520 1.680 17.360 1.960 ;
      LAYER met1 ;
        RECT 17.360 1.680 18.760 1.960 ;
        RECT 0.000 0.560 2.240 1.680 ;
      LAYER met1 ;
        RECT 2.240 1.400 16.800 1.680 ;
      LAYER met1 ;
        RECT 16.800 1.400 18.760 1.680 ;
      LAYER met1 ;
        RECT 2.240 1.120 15.680 1.400 ;
      LAYER met1 ;
        RECT 15.680 1.120 18.760 1.400 ;
      LAYER met1 ;
        RECT 2.240 0.840 14.560 1.120 ;
      LAYER met1 ;
        RECT 14.560 0.840 18.760 1.120 ;
      LAYER met1 ;
        RECT 2.240 0.560 14.280 0.840 ;
      LAYER met1 ;
        RECT 14.280 0.560 18.760 0.840 ;
        RECT 0.000 0.280 2.520 0.560 ;
      LAYER met1 ;
        RECT 2.520 0.280 14.000 0.560 ;
      LAYER met1 ;
        RECT 14.000 0.280 18.760 0.560 ;
        RECT 0.000 0.000 6.160 0.280 ;
      LAYER met1 ;
        RECT 6.160 0.000 13.440 0.280 ;
      LAYER met1 ;
        RECT 13.440 0.000 18.760 0.280 ;
      LAYER met2 ;
        RECT 0.000 27.440 7.560 27.720 ;
      LAYER met2 ;
        RECT 7.560 27.440 8.120 27.720 ;
      LAYER met2 ;
        RECT 0.000 27.160 7.000 27.440 ;
      LAYER met2 ;
        RECT 7.000 27.160 8.120 27.440 ;
      LAYER met2 ;
        RECT 0.000 26.880 6.720 27.160 ;
      LAYER met2 ;
        RECT 6.720 26.880 8.120 27.160 ;
      LAYER met2 ;
        RECT 0.000 26.600 6.440 26.880 ;
      LAYER met2 ;
        RECT 6.440 26.600 8.120 26.880 ;
      LAYER met2 ;
        RECT 0.000 26.320 6.160 26.600 ;
      LAYER met2 ;
        RECT 6.160 26.320 8.120 26.600 ;
      LAYER met2 ;
        RECT 0.000 26.040 5.880 26.320 ;
      LAYER met2 ;
        RECT 5.880 26.040 8.120 26.320 ;
      LAYER met2 ;
        RECT 8.120 26.040 18.760 27.720 ;
        RECT 0.000 25.480 5.600 26.040 ;
      LAYER met2 ;
        RECT 5.600 25.480 8.120 26.040 ;
      LAYER met2 ;
        RECT 8.120 25.760 11.480 26.040 ;
      LAYER met2 ;
        RECT 11.480 25.760 12.040 26.040 ;
      LAYER met2 ;
        RECT 8.120 25.480 10.920 25.760 ;
      LAYER met2 ;
        RECT 10.920 25.480 12.040 25.760 ;
      LAYER met2 ;
        RECT 0.000 24.920 5.320 25.480 ;
      LAYER met2 ;
        RECT 5.320 24.920 7.840 25.480 ;
      LAYER met2 ;
        RECT 7.840 25.200 10.080 25.480 ;
      LAYER met2 ;
        RECT 10.080 25.200 12.040 25.480 ;
      LAYER met2 ;
        RECT 7.840 24.920 9.800 25.200 ;
      LAYER met2 ;
        RECT 9.800 24.920 12.040 25.200 ;
      LAYER met2 ;
        RECT 12.040 24.920 18.760 26.040 ;
        RECT 0.000 24.080 5.040 24.920 ;
      LAYER met2 ;
        RECT 5.040 24.640 7.840 24.920 ;
      LAYER met2 ;
        RECT 7.840 24.640 9.240 24.920 ;
      LAYER met2 ;
        RECT 9.240 24.640 11.760 24.920 ;
        RECT 5.040 24.080 7.560 24.640 ;
      LAYER met2 ;
        RECT 7.560 24.360 8.960 24.640 ;
      LAYER met2 ;
        RECT 8.960 24.360 11.760 24.640 ;
      LAYER met2 ;
        RECT 7.560 24.080 8.400 24.360 ;
      LAYER met2 ;
        RECT 8.400 24.080 11.760 24.360 ;
      LAYER met2 ;
        RECT 11.760 24.080 18.760 24.920 ;
        RECT 0.000 21.560 4.760 24.080 ;
      LAYER met2 ;
        RECT 4.760 23.800 7.560 24.080 ;
      LAYER met2 ;
        RECT 7.560 23.800 8.120 24.080 ;
      LAYER met2 ;
        RECT 8.120 23.800 11.480 24.080 ;
        RECT 4.760 23.240 7.280 23.800 ;
      LAYER met2 ;
        RECT 7.280 23.520 7.840 23.800 ;
      LAYER met2 ;
        RECT 7.840 23.520 11.480 23.800 ;
      LAYER met2 ;
        RECT 11.480 23.520 18.760 24.080 ;
        RECT 7.280 23.240 7.560 23.520 ;
      LAYER met2 ;
        RECT 7.560 23.240 11.200 23.520 ;
        RECT 4.760 22.960 11.200 23.240 ;
      LAYER met2 ;
        RECT 11.200 22.960 18.760 23.520 ;
      LAYER met2 ;
        RECT 4.760 22.680 10.920 22.960 ;
      LAYER met2 ;
        RECT 10.920 22.680 18.760 22.960 ;
      LAYER met2 ;
        RECT 4.760 22.120 10.640 22.680 ;
      LAYER met2 ;
        RECT 10.640 22.120 18.760 22.680 ;
      LAYER met2 ;
        RECT 4.760 21.840 10.360 22.120 ;
      LAYER met2 ;
        RECT 10.360 21.840 18.760 22.120 ;
      LAYER met2 ;
        RECT 4.760 21.560 10.080 21.840 ;
      LAYER met2 ;
        RECT 10.080 21.560 18.760 21.840 ;
        RECT 0.000 21.280 3.920 21.560 ;
      LAYER met2 ;
        RECT 3.920 21.280 9.800 21.560 ;
      LAYER met2 ;
        RECT 9.800 21.280 18.760 21.560 ;
        RECT 0.000 21.000 3.080 21.280 ;
      LAYER met2 ;
        RECT 3.080 21.000 9.520 21.280 ;
      LAYER met2 ;
        RECT 9.520 21.000 18.760 21.280 ;
        RECT 0.000 20.720 2.800 21.000 ;
      LAYER met2 ;
        RECT 2.800 20.720 8.960 21.000 ;
      LAYER met2 ;
        RECT 8.960 20.720 18.760 21.000 ;
        RECT 0.000 20.440 2.240 20.720 ;
      LAYER met2 ;
        RECT 2.240 20.440 8.680 20.720 ;
      LAYER met2 ;
        RECT 8.680 20.440 18.760 20.720 ;
        RECT 0.000 20.160 1.960 20.440 ;
      LAYER met2 ;
        RECT 1.960 20.160 8.120 20.440 ;
      LAYER met2 ;
        RECT 0.000 19.880 1.680 20.160 ;
      LAYER met2 ;
        RECT 1.680 19.880 8.120 20.160 ;
      LAYER met2 ;
        RECT 0.000 19.600 1.400 19.880 ;
      LAYER met2 ;
        RECT 1.400 19.600 8.120 19.880 ;
      LAYER met2 ;
        RECT 8.120 19.600 18.760 20.440 ;
        RECT 0.000 19.320 1.120 19.600 ;
      LAYER met2 ;
        RECT 1.120 19.320 8.400 19.600 ;
      LAYER met2 ;
        RECT 0.000 19.040 0.840 19.320 ;
      LAYER met2 ;
        RECT 0.840 19.040 8.400 19.320 ;
      LAYER met2 ;
        RECT 0.000 18.760 0.560 19.040 ;
      LAYER met2 ;
        RECT 0.560 18.760 8.400 19.040 ;
      LAYER met2 ;
        RECT 0.000 18.480 0.280 18.760 ;
      LAYER met2 ;
        RECT 0.280 18.480 8.400 18.760 ;
        RECT 0.000 17.360 8.400 18.480 ;
      LAYER met2 ;
        RECT 0.000 16.800 0.280 17.360 ;
      LAYER met2 ;
        RECT 0.280 16.800 8.400 17.360 ;
      LAYER met2 ;
        RECT 8.400 16.800 18.760 19.600 ;
        RECT 0.000 16.240 0.560 16.800 ;
      LAYER met2 ;
        RECT 0.560 16.520 8.680 16.800 ;
      LAYER met2 ;
        RECT 8.680 16.520 18.760 16.800 ;
      LAYER met2 ;
        RECT 0.560 16.240 9.240 16.520 ;
      LAYER met2 ;
        RECT 9.240 16.240 18.760 16.520 ;
        RECT 0.000 15.960 0.840 16.240 ;
      LAYER met2 ;
        RECT 0.840 15.960 9.800 16.240 ;
      LAYER met2 ;
        RECT 9.800 15.960 18.760 16.240 ;
        RECT 0.000 15.680 1.400 15.960 ;
      LAYER met2 ;
        RECT 1.400 15.680 10.360 15.960 ;
      LAYER met2 ;
        RECT 10.360 15.680 18.760 15.960 ;
        RECT 0.000 14.280 2.520 15.680 ;
      LAYER met2 ;
        RECT 2.520 15.400 10.920 15.680 ;
      LAYER met2 ;
        RECT 10.920 15.400 18.760 15.680 ;
      LAYER met2 ;
        RECT 2.520 15.120 11.200 15.400 ;
      LAYER met2 ;
        RECT 11.200 15.120 18.760 15.400 ;
      LAYER met2 ;
        RECT 2.520 14.840 11.760 15.120 ;
      LAYER met2 ;
        RECT 11.760 14.840 18.760 15.120 ;
      LAYER met2 ;
        RECT 2.520 14.560 12.040 14.840 ;
      LAYER met2 ;
        RECT 12.040 14.560 18.760 14.840 ;
      LAYER met2 ;
        RECT 2.520 14.280 12.600 14.560 ;
      LAYER met2 ;
        RECT 12.600 14.280 18.760 14.560 ;
        RECT 0.000 9.240 2.240 14.280 ;
      LAYER met2 ;
        RECT 2.240 14.000 12.880 14.280 ;
      LAYER met2 ;
        RECT 12.880 14.000 18.760 14.280 ;
      LAYER met2 ;
        RECT 2.240 13.720 13.160 14.000 ;
      LAYER met2 ;
        RECT 13.160 13.720 18.760 14.000 ;
      LAYER met2 ;
        RECT 2.240 13.440 13.440 13.720 ;
      LAYER met2 ;
        RECT 13.440 13.440 18.760 13.720 ;
      LAYER met2 ;
        RECT 2.240 13.160 13.720 13.440 ;
      LAYER met2 ;
        RECT 13.720 13.160 18.760 13.440 ;
      LAYER met2 ;
        RECT 2.240 12.880 14.000 13.160 ;
      LAYER met2 ;
        RECT 14.000 12.880 18.760 13.160 ;
      LAYER met2 ;
        RECT 2.240 12.600 14.280 12.880 ;
      LAYER met2 ;
        RECT 14.280 12.600 18.760 12.880 ;
      LAYER met2 ;
        RECT 2.240 12.320 14.560 12.600 ;
      LAYER met2 ;
        RECT 14.560 12.320 18.760 12.600 ;
      LAYER met2 ;
        RECT 2.240 12.040 14.840 12.320 ;
      LAYER met2 ;
        RECT 14.840 12.040 18.760 12.320 ;
      LAYER met2 ;
        RECT 2.240 11.760 15.120 12.040 ;
      LAYER met2 ;
        RECT 15.120 11.760 18.760 12.040 ;
      LAYER met2 ;
        RECT 2.240 11.480 15.400 11.760 ;
      LAYER met2 ;
        RECT 15.400 11.480 18.760 11.760 ;
      LAYER met2 ;
        RECT 2.240 11.200 15.680 11.480 ;
      LAYER met2 ;
        RECT 15.680 11.200 18.760 11.480 ;
      LAYER met2 ;
        RECT 2.240 10.640 15.960 11.200 ;
      LAYER met2 ;
        RECT 15.960 10.640 18.760 11.200 ;
      LAYER met2 ;
        RECT 2.240 10.360 16.240 10.640 ;
      LAYER met2 ;
        RECT 16.240 10.360 18.760 10.640 ;
      LAYER met2 ;
        RECT 2.240 9.800 16.520 10.360 ;
      LAYER met2 ;
        RECT 16.520 9.800 18.760 10.360 ;
      LAYER met2 ;
        RECT 2.240 9.240 16.800 9.800 ;
      LAYER met2 ;
        RECT 16.800 9.240 18.760 9.800 ;
        RECT 0.000 8.400 2.520 9.240 ;
      LAYER met2 ;
        RECT 2.520 8.680 17.080 9.240 ;
      LAYER met2 ;
        RECT 17.080 8.680 18.760 9.240 ;
      LAYER met2 ;
        RECT 2.520 8.400 17.360 8.680 ;
      LAYER met2 ;
        RECT 0.000 7.840 2.800 8.400 ;
      LAYER met2 ;
        RECT 2.800 8.120 17.360 8.400 ;
      LAYER met2 ;
        RECT 17.360 8.120 18.760 8.680 ;
      LAYER met2 ;
        RECT 2.800 7.840 17.640 8.120 ;
      LAYER met2 ;
        RECT 0.000 3.920 3.360 7.840 ;
      LAYER met2 ;
        RECT 3.360 7.000 17.640 7.840 ;
      LAYER met2 ;
        RECT 17.640 7.000 18.760 8.120 ;
      LAYER met2 ;
        RECT 3.360 4.200 17.920 7.000 ;
      LAYER met2 ;
        RECT 17.920 4.200 18.760 7.000 ;
      LAYER met2 ;
        RECT 3.360 3.920 18.480 4.200 ;
      LAYER met2 ;
        RECT 18.480 3.920 18.760 4.200 ;
        RECT 0.000 2.240 3.640 3.920 ;
      LAYER met2 ;
        RECT 3.640 3.080 18.760 3.920 ;
        RECT 3.640 2.800 18.480 3.080 ;
      LAYER met2 ;
        RECT 18.480 2.800 18.760 3.080 ;
      LAYER met2 ;
        RECT 3.640 2.240 17.920 2.800 ;
      LAYER met2 ;
        RECT 17.920 2.240 18.760 2.800 ;
        RECT 0.000 1.960 2.800 2.240 ;
      LAYER met2 ;
        RECT 2.800 1.960 17.640 2.240 ;
      LAYER met2 ;
        RECT 17.640 1.960 18.760 2.240 ;
        RECT 0.000 1.680 2.520 1.960 ;
      LAYER met2 ;
        RECT 2.520 1.680 17.360 1.960 ;
      LAYER met2 ;
        RECT 17.360 1.680 18.760 1.960 ;
        RECT 0.000 0.560 2.240 1.680 ;
      LAYER met2 ;
        RECT 2.240 1.400 16.800 1.680 ;
      LAYER met2 ;
        RECT 16.800 1.400 18.760 1.680 ;
      LAYER met2 ;
        RECT 2.240 1.120 15.680 1.400 ;
      LAYER met2 ;
        RECT 15.680 1.120 18.760 1.400 ;
      LAYER met2 ;
        RECT 2.240 0.840 14.560 1.120 ;
      LAYER met2 ;
        RECT 14.560 0.840 18.760 1.120 ;
      LAYER met2 ;
        RECT 2.240 0.560 14.280 0.840 ;
      LAYER met2 ;
        RECT 14.280 0.560 18.760 0.840 ;
        RECT 0.000 0.280 2.520 0.560 ;
      LAYER met2 ;
        RECT 2.520 0.280 14.000 0.560 ;
      LAYER met2 ;
        RECT 14.000 0.280 18.760 0.560 ;
        RECT 0.000 0.000 6.160 0.280 ;
      LAYER met2 ;
        RECT 6.160 0.000 13.440 0.280 ;
      LAYER met2 ;
        RECT 13.440 0.000 18.760 0.280 ;
      LAYER met3 ;
        RECT 0.000 0.000 18.760 27.720 ;
      LAYER met4 ;
        RECT 0.000 0.000 18.760 27.720 ;
      LAYER met5 ;
        RECT 0.000 0.000 18.760 27.720 ;
  END
END white_rabbit
END LIBRARY

